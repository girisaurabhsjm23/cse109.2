* C:\Users\User\Documents\Schematic4.sch

* Schematics Version 9.1 - Web Update 1
* Thu Aug 17 10:48:49 2023



** Analysis setup **
.ac DEC 10 0.1 1gig
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic4.net"
.INC "Schematic4.als"


.probe


.END

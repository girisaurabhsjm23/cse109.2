* C:\Users\User\Documents\Schematic2.sch

* Schematics Version 9.1 - Web Update 1
* Thu Aug 10 11:02:50 2023



** Analysis setup **
.tran 0ns 100ms
.OP 


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "Schematic2.net"
.INC "Schematic2.als"


.probe


.END
